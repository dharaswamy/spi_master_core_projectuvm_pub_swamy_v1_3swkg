
`define NO_SLAVES 8 
`define WB_ADDR_WIDTH 5


//nagesh sir 2 months
//sastri sir    8 months
